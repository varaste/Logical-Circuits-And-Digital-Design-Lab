module bcd_to_gray(a, b);
input [3:0]  a;
output [3:0] b;

and #10 (b[3], a[3],a[3]);
xor #10 (b[2],a[3],a[2]);
xor #10 (b[1], a[2],a[1]);
xor #10 (b[0], a[1], a[0]);
endmodule



module gray_to_bcd(a, b);
input [3:0]  a;
output [3:0] b;

and #10 (b[3], a[3],a[3]);
xor #10 (b[2],b[3],a[2]);
xor #10 (b[1], b[2],a[1]);
xor #10 (b[0], b[1], a[0]);
endmodule




module test_cicuit;
reg [3:0] a;
wire[3:0] b;


gray_to_bcd bin(a,b);
initial
begin
a[3]=1'b0; a[2]=1'b0; a[1]=1'b0; a[0]=1'b0;
#100
a[3]=1'b0; a[2]=1'b0; a[1]=1'b0; a[0]=1'b1;
#100
a[3]=1'b0; a[2]=1'b0; a[1]=1'b1; a[0]=1'b0;
#100
a[3]=1'b0; a[2]=1'b0; a[1]=1'b1; a[0]=1'b1;
#100
a[3]=1'b0; a[2]=1'b1; a[1]=1'b0; a[0]=1'b0;
#100
a[3]=1'b0; a[2]=1'b1; a[1]=1'b0; a[0]=1'b1;
#100
a[3]=1'b0; a[2]=1'b1; a[1]=1'b1; a[0]=1'b0;
#100
a[3]=1'b0; a[2]=1'b1; a[1]=1'b1; a[0]=1'b1;
#100
a[3]=1'b1; a[2]=1'b0; a[1]=1'b0; a[0]=1'b0;
#100
a[3]=1'b1; a[2]=1'b0; a[1]=1'b0; a[0]=1'b1;
#100
a[3]=1'b1; a[2]=1'b0; a[1]=1'b1; a[0]=1'b0;
#100
a[3]=1'b1; a[2]=1'b0; a[1]=1'b1; a[0]=1'b1;
#100
a[3]=1'b1; a[2]=1'b1; a[1]=1'b0; a[0]=1'b0;
#100
a[3]=1'b1; a[2]=1'b1; a[1]=1'b0; a[0]=1'b1;
#100
a[3]=1'b1; a[2]=1'b1; a[1]=1'b1; a[0]=1'b0;
#100
a[3]=1'b1; a[2]=1'b1; a[1]=1'b1; a[0]=1'b1;
#100
$finish;

end
endmodule


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:08:33 11/21/2017 
// Design Na//////////////////////////////////////////////////////////////////////////////////
module uut(
    );


endmodule
